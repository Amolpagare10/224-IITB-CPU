library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity shifter_1_bit is 
	port (input: in std_logic_vector(15 downto 0);
			alu_b: out std_logic_vector(15 downto 0);
			s: in std_logic_vector(3 downto 0);
			clk: in std_logic
	);
	end entity;
	
architecture exe of shifter_1_bit is
begin
	lshift_1_bit_proc: process(input,s, clk)
	variable i: integer;
	begin
	 if (s="1100") then
	 alu_b(0) <= '0';
		 FOR i IN 0 TO 14 LOOP
	        alu_b(i+1) <= input(i);
	      END LOOP;
	end if;
	end process;
end exe;